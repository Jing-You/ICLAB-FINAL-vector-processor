module MEM_stage();
endmodule
