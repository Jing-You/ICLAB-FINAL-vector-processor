module WB_stage();

endmodule