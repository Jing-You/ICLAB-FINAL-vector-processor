module MEM_WB_stage();

endmodule;